module pwm #(
    parameters
) (
   input ; 
);
    
endmodule